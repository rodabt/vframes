module vframes
